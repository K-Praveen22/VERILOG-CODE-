module arithmatic_op;
  reg[3:0]i1,i2;
  initial begin
    i1=4'h6;
    i2=4'h2;
    $display("i1=%0h and i2=%0h",i1,i2);
    $display("add:%0h",i1+i2);
    $display("sub;%0h",i1-i2);
    $display("mul:%0h",i1*i2);
    $display("div:%0h",i1/i2);
    $display("pow:%0h",i1**3);
    $display("mod:%0h",i1%i2);
    
    i1=4'ha; i2=4'h3;
    
    $display("\nil=%0h and i2=%oh",i1,i2);
    $display("mod:%0h",i1,i2);
  end
endmodule  
